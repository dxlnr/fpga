module baud_rate_generator_tb();
endmodule
